library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL;

ENTITY regbank IS
	PORT(
			INSTR2,INSTR3, INSTRD : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			WRITEFLAG: IN STD_LOGIC;
			WRITEBACKDATA: IN STD_LOGIC_VECTOR(15 DOWNTO 0);
			OUTREG1,OUTREG2 : OUT STD_LOGIC_VECTOR(15 DOWNTO 0)
	);
END regbank;

ARCHITECTURE behavior OF regbank IS

	TYPE BANK IS ARRAY(0 TO 15) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL BANKREG : BANK;
	
		BEGIN 
			OUTREG1 <= BANKREG( TO_INTEGER(UNSIGNED(INSTR2)));
			OUTREG2 <= BANKREG( TO_INTEGER(UNSIGNED(INSTR3)));
			PROCESS(WRITEFLAG)
				BEGIN
					IF WRITEFLAG = '1' THEN
						BANKREG(TO_INTEGER( UNSIGNED(INSTRD))) <= WRITEBACKDATA;
					END IF;
			END PROCESS;
			
END behavior;